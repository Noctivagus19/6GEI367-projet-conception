LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_UNSIGNED.ALL; 


ENTITY psa IS
	PORT (D0, D1 : IN STD_LOGIC;
			SEL : IN STD_LOGIC;
			MX_OUT : OUT STD_LOGIC);
END psa;

ARCHITECTURE rtl OF psa IS
BEGIN
	WITH SEL select
		MX_OUT <= D0 WHEN '0',
				D1 WHEN '1',
				'0' WHEN OTHERS;
END rtl;